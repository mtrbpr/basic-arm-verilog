module instruction_memory(
    input [31:0] addr,
    input rst,
    output [31:0] instruction
);

reg [31:0] mem [0:1023];

always @(rst) begin
    mem[0] <= 32'b11100011101000000000000000010100;
    mem[1] <= 32'b11100011101000000001101000000001;
    mem[2] <= 32'b11100011101000000010000100000011;
    mem[3] <= 32'b11100000100100100011000000000010;
    mem[4] <= 32'b11100000101000000100000000000000;
    mem[5] <= 32'b11100000010001000101000100000100;
    mem[6] <= 32'b11100000110000000110000010100000;
    mem[7] <= 32'b11100001100001010111000101000010;
    mem[8] <= 32'b11100000000001111000000000000011;
    mem[9] <= 32'b11100001111000001001000000000110;
    mem[10] <= 32'b11100000001001001010000000000101;
    mem[11] <= 32'b11100001010110000000000000000110;
    mem[12] <= 32'b00010000100000010001000000000001;
    mem[13] <= 32'b11100001000110010000000000001000;
    mem[14] <= 32'b00000000100000100010000000000010;
    mem[15] <= 32'b11100011101000000000101100000001;
    mem[16] <= 32'b11100100100000000001000000000000;
    mem[17] <= 32'b11100100100100001011000000000000;
    mem[18] <= 32'b11100100100000000010000000000100;
    mem[19] <= 32'b11100100100000000011000000001000;
    mem[20] <= 32'b11100100100000000100000000001101;
    mem[21] <= 32'b11100100100000000101000000010000;
    mem[22] <= 32'b11100100100000000110000000010100;
    mem[23] <= 32'b11100100100100001010000000000100;
    mem[24] <= 32'b11100100100000000111000000011000;
    mem[25] <= 32'b11100011101000000001000000000100;
    mem[26] <= 32'b11100011101000000010000000000000;
    mem[27] <= 32'b11100011101000000011000000000000;
    mem[28] <= 32'b11100000100000000100000100000011;
    mem[29] <= 32'b11100100100101000101000000000000;
    mem[30] <= 32'b11100100100101000110000000000100;
    mem[31] <= 32'b11100001010101010000000000000110;
    mem[32] <= 32'b11000100100001000110000000000000;
    mem[33] <= 32'b11000100100001000101000000000100;
    mem[34] <= 32'b11100010100000110011000000000001;
    mem[35] <= 32'b11100011010100110000000000000011;
    mem[36] <= 32'b10111010111111111111111111110111;
    mem[37] <= 32'b11100010100000100010000000000001;
    mem[38] <= 32'b11100001010100100000000000000001;
    mem[39] <= 32'b10111010111111111111111111110011;
    mem[40] <= 32'b11100100100100000001000000000000;
    mem[41] <= 32'b11100100100100000010000000000100;
    mem[42] <= 32'b11100100100100000011000000001000;
    mem[43] <= 32'b11100100100100000100000000001100;
    mem[44] <= 32'b11100100100100000101000000010000;
    mem[45] <= 32'b11100100100100000110000000010100;
    mem[46] <= 32'b11101010111111111111111111111111;
end

/*initial begin
    $readmemb("./instruction_fetch/instructions.txt", mem);
end*/
assign instruction = rst ? 32'b0 : mem[addr >> 2];

endmodule